library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity SLL2 is 
	generic(
		width : positive := 32
	);
	port(
		in0	: in std_logic_vector(width-1 downto 0);
		out0 : out std_logic_vector(width-1 downto 0)
	);
end SLL2;

architecture BHV of SLL2 is
begin
	out0 <= std_logic_vector(unsigned(in0) sll 2);
end BHV; 
